package dst_agent_main;

endpackage

